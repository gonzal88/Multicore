mg221@cparch03.ecn.purdue.edu.13699:1447956357