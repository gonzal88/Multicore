mg221@cparch07.ecn.purdue.edu.9255:1441056760