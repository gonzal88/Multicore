mg221@cparch04.ecn.purdue.edu.6452:1446132498