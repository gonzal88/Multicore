mg221@cparch16.ecn.purdue.edu.5751:1445381375